`timescale 1ns/1ps

module forwarding_unit(
    input [2:0] id_ex_rs1,
    input [2:0] id_ex_rs2,
    input [2:0] ex_mem_rd,
    input [2:0] mem_wb_rd,
    input ex_mem_regwrite,
    input mem_wb_regwrite,
    output reg [1:0] forwardA,
    output reg [1:0] forwardB
);
    always @* begin
        forwardA = 2'b00;
        forwardB = 2'b00;
        if (ex_mem_regwrite && (ex_mem_rd != 3'b000) && (ex_mem_rd == id_ex_rs1))
            forwardA = 2'b01;
        if (ex_mem_regwrite && (ex_mem_rd != 3'b000) && (ex_mem_rd == id_ex_rs2))
            forwardB = 2'b01;
        if (mem_wb_regwrite && (mem_wb_rd != 3'b000) && (mem_wb_rd == id_ex_rs1) &&
            !(ex_mem_regwrite && (ex_mem_rd != 3'b000) && (ex_mem_rd == id_ex_rs1)))
            forwardA = 2'b10;
        if (mem_wb_regwrite && (mem_wb_rd != 3'b000) && (mem_wb_rd == id_ex_rs2) &&
            !(ex_mem_regwrite && (ex_mem_rd != 3'b000) && (ex_mem_rd == id_ex_rs2)))
            forwardB = 2'b10;
    end
endmodule
